module logic1(
    output logic Q
);
    assign Q = 1'b1;
endmodule