module logic0(
    output logic Q
);
    assign Q = 1'b0;
endmodule